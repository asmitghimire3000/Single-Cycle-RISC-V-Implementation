// module PC_target_calc(PC1,PC2,PCT);
//     input [31:0] PC1;
//     input [31:0] PC2;
//     output [31:0] PCT;

//     assign PCT = PC1 + PC2;
// endmodule